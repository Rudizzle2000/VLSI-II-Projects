
module gcd_clk_gen_ds 
    (
      input reset_i,          // Reset signal for the GCD module
      input clk_reset_i,      // Reset signal for the clock generator module
      input ds_reset_i,       // Reset signal for the data source module
      input [7:0] select_i,   // Configuration input to select clock generation parameters

      input [63:0] data_i,    // Input data to the GCD module
      input v_i,              // Valid signal indicating that input data is valid
      output ready_o,         // Output signal indicating that the GCD module is ready to accept data
      output clk_o,           // Output clock signal generated by the clock generator module

      output logic [63:0] data_o, // Output data from the GCD module
      output logic v_o,           // Valid signal indicating that the output data is valid
      input yumi_i                // Yumi signal for handshaking with the GCD module
    );

    // Instantiate the clock generator and data source module (clk_gen_ds)
    // This module generates the clock signal based on the reset signals and
    // the select input.
    clk_gen_ds 
    CGDS (
          .clk_reset_i(clk_reset_i),  // Clock generator reset input
          .ds_reset_i(ds_reset_i),    // Data source reset input
          .select_i(select_i),        // Clock generation configuration input
          .clk_o(clk_o),              // Clock output generated by the module
          .ds_enable()                // Data source enable signal (ignored in this case, used only for waveform observation)
    );

    // Instantiate the GCD module
    // This module computes the greatest common divisor (GCD) of the input data.
    gcd
    GCD (
         .clk_i(clk_o),            // Clock input to the GCD module
         .reset_i(reset_i),        // Reset input to the GCD module
         .data_in(data_i),         // Input data to the GCD module
         .v_i(v_i),                // Valid signal indicating input data is valid
         .ready_o(ready_o),        // Output signal indicating that GCD is ready to accept data
         .data_out(data_o),        // Output data from the GCD module
         .v_o(v_o),                // Valid signal indicating output data is valid
         .yumi_i(yumi_i)           // Yumi signal for handshaking with the GCD module
    );

endmodule
